library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package neorv32_dcache_memory_tb_pkg is

	constant cache_size : integer := 512;

	type ext_mem_type is array (0 to 1023) of std_ulogic_vector(31 downto 0);

	constant cache_ext_mem : ext_mem_type := (
		00000000 => x"06b3d9b3",
		00000001 => x"22433ed9",
		00000002 => x"0b28eed7",
		00000003 => x"626d29be",
		00000004 => x"34207f83",
		00000005 => x"221e6f79",
		00000006 => x"0dc91f05",
		00000007 => x"6b54154a",
		00000008 => x"735a7c19",
		00000009 => x"6ffa4a47",
		00000010 => x"04e2382a",
		00000011 => x"3087256a",
		00000012 => x"44a244be",
		00000013 => x"47fa0f46",
		00000014 => x"2a857444",
		00000015 => x"2b9f46bb",
		00000016 => x"6d112ca7",
		00000017 => x"06a4b6a5",
		00000018 => x"146fd14c",
		00000019 => x"11499016",
		00000020 => x"2b29ea5e",
		00000021 => x"47cd9a64",
		00000022 => x"2ab9d716",
		00000023 => x"59d0f898",
		00000024 => x"1f618346",
		00000025 => x"14f6a3ce",
		00000026 => x"0036bd9a",
		00000027 => x"73f4b6aa",
		00000028 => x"37d7e290",
		00000029 => x"6304ee5d",
		00000030 => x"0b36eb41",
		00000031 => x"7076f578",
		00000032 => x"4c7e23a1",
		00000033 => x"30550698",
		00000034 => x"08f1ba77",
		00000035 => x"00d81b37",
		00000036 => x"2860f5a2",
		00000037 => x"5db37659",
		00000038 => x"39629b19",
		00000039 => x"0d0f8a0d",
		00000040 => x"73e41a69",
		00000041 => x"059e1aa6",
		00000042 => x"0bdfb58c",
		00000043 => x"5564c896",
		00000044 => x"1232caef",
		00000045 => x"1028f338",
		00000046 => x"652112fb",
		00000047 => x"740bbaf9",
		00000048 => x"02b7dc42",
		00000049 => x"2559c082",
		00000050 => x"74a094ca",
		00000051 => x"371f21e1",
		00000052 => x"49656fa8",
		00000053 => x"3d0bd352",
		00000054 => x"21f60fc2",
		00000055 => x"3c11c846",
		00000056 => x"6b3e4390",
		00000057 => x"04b4017b",
		00000058 => x"6267ddc5",
		00000059 => x"270d6c3f",
		00000060 => x"2bf69168",
		00000061 => x"42c61737",
		00000062 => x"669770b1",
		00000063 => x"3dd1acba",
		00000064 => x"1a7a7820",
		00000065 => x"691f71e4",
		00000066 => x"4df08497",
		00000067 => x"51c2c66f",
		00000068 => x"43773120",
		00000069 => x"484bd381",
		00000070 => x"67986796",
		00000071 => x"7af3bea6",
		00000072 => x"285a8b02",
		00000073 => x"019b2d04",
		00000074 => x"32f977bb",
		00000075 => x"724be697",
		00000076 => x"6277bcbc",
		00000077 => x"52b53161",
		00000078 => x"41a1dca3",
		00000079 => x"3799fb84",
		00000080 => x"57a8bef8",
		00000081 => x"44ee3467",
		00000082 => x"51b58f43",
		00000083 => x"65f2a614",
		00000084 => x"55550988",
		00000085 => x"4c5a42ef",
		00000086 => x"71eebffd",
		00000087 => x"6ab07b25",
		00000088 => x"3e39b846",
		00000089 => x"42a350d4",
		00000090 => x"55906ea4",
		00000091 => x"35b20d9d",
		00000092 => x"2ff0532c",
		00000093 => x"4149d990",
		00000094 => x"04136034",
		00000095 => x"6c75b209",
		00000096 => x"6088bf17",
		00000097 => x"529e2663",
		00000098 => x"173a3e0f",
		00000099 => x"5ce7ed32",
		00000100 => x"68fbfdf2",
		00000101 => x"0a92f4e9",
		00000102 => x"74f2596e",
		00000103 => x"3e52e876",
		00000104 => x"543bc629",
		00000105 => x"21858582",
		00000106 => x"15c6b7c0",
		00000107 => x"2ade0534",
		00000108 => x"2b201187",
		00000109 => x"46f0254f",
		00000110 => x"32129f41",
		00000111 => x"71242ddb",
		00000112 => x"0961979b",
		00000113 => x"5c8efa32",
		00000114 => x"3a7757ec",
		00000115 => x"319eb312",
		00000116 => x"495d95fe",
		00000117 => x"63adb498",
		00000118 => x"2b05865c",
		00000119 => x"021663e1",
		00000120 => x"18332de1",
		00000121 => x"4b08a8b6",
		00000122 => x"0b48bcf1",
		00000123 => x"6a71fed2",
		00000124 => x"506cb56f",
		00000125 => x"2e87abc0",
		00000126 => x"01a4625e",
		00000127 => x"72b50758",
		00000128 => x"2d0b81e2",
		00000129 => x"7fafcd7b",
		00000130 => x"1d541fc6",
		00000131 => x"33ee986b",
		00000132 => x"44187e63",
		00000133 => x"4021049b",
		00000134 => x"5ca10027",
		00000135 => x"697bcf17",
		00000136 => x"745f2279",
		00000137 => x"07a51c73",
		00000138 => x"51c439d8",
		00000139 => x"24d36df6",
		00000140 => x"7ef31381",
		00000141 => x"3f54ef29",
		00000142 => x"7b664a72",
		00000143 => x"61d0e5de",
		00000144 => x"50a3891d",
		00000145 => x"5c32a6d9",
		00000146 => x"1ddf2c25",
		00000147 => x"45a75dbf",
		00000148 => x"3ded88da",
		00000149 => x"7d86beb2",
		00000150 => x"16bb42ac",
		00000151 => x"13ae766e",
		00000152 => x"7ef878ef",
		00000153 => x"44a819b9",
		00000154 => x"38e55f98",
		00000155 => x"3075a47b",
		00000156 => x"60361287",
		00000157 => x"3b0bbfd4",
		00000158 => x"05a60c1b",
		00000159 => x"014ca9b5",
		00000160 => x"113ec10c",
		00000161 => x"3a695c14",
		00000162 => x"18ba05e9",
		00000163 => x"02b06a70",
		00000164 => x"20d07b32",
		00000165 => x"6641fda3",
		00000166 => x"2d0fe4bb",
		00000167 => x"57acfa50",
		00000168 => x"22ce98e2",
		00000169 => x"7a32b220",
		00000170 => x"37961ced",
		00000171 => x"512fb538",
		00000172 => x"35ce44c5",
		00000173 => x"000ba4c3",
		00000174 => x"0de74998",
		00000175 => x"4f0d0367",
		00000176 => x"0803907b",
		00000177 => x"41522ccc",
		00000178 => x"2d72a741",
		00000179 => x"5a80b275",
		00000180 => x"0b5d6f56",
		00000181 => x"0a9ca5df",
		00000182 => x"37731b96",
		00000183 => x"72e09b41",
		00000184 => x"011888a2",
		00000185 => x"65daa143",
		00000186 => x"449520b9",
		00000187 => x"30509219",
		00000188 => x"0967ec61",
		00000189 => x"45f66db7",
		00000190 => x"58dbbd49",
		00000191 => x"514abb48",
		00000192 => x"33bd1053",
		00000193 => x"03bac1c0",
		00000194 => x"7e1fe39e",
		00000195 => x"29464d73",
		00000196 => x"219ae945",
		00000197 => x"7a568b15",
		00000198 => x"3c7b3b6f",
		00000199 => x"043a5d63",
		00000200 => x"601ab435",
		00000201 => x"47e21f64",
		00000202 => x"2adbba2f",
		00000203 => x"35004c31",
		00000204 => x"2c974a62",
		00000205 => x"030b9fe9",
		00000206 => x"51cef1be",
		00000207 => x"516b32a6",
		00000208 => x"7c1eac61",
		00000209 => x"14f9517d",
		00000210 => x"7122fbf9",
		00000211 => x"7b497f8d",
		00000212 => x"35a3080a",
		00000213 => x"08393ab8",
		00000214 => x"5bde2e28",
		00000215 => x"6f5308c3",
		00000216 => x"56eb2caa",
		00000217 => x"126e12d2",
		00000218 => x"2fa149bf",
		00000219 => x"5599f486",
		00000220 => x"1e134823",
		00000221 => x"5f3f20ba",
		00000222 => x"0a083d83",
		00000223 => x"6991a28c",
		00000224 => x"70801689",
		00000225 => x"5052a569",
		00000226 => x"0750fe30",
		00000227 => x"610834c7",
		00000228 => x"4264a27e",
		00000229 => x"31900d0a",
		00000230 => x"44cdfdfe",
		00000231 => x"27305fcd",
		00000232 => x"12b4b0b8",
		00000233 => x"74f4d8b6",
		00000234 => x"53f59203",
		00000235 => x"62dfb063",
		00000236 => x"7539b1c2",
		00000237 => x"2545dfaa",
		00000238 => x"6358533a",
		00000239 => x"6af76489",
		00000240 => x"31d33f68",
		00000241 => x"2f2a9eff",
		00000242 => x"10302ae0",
		00000243 => x"447846c9",
		00000244 => x"7cca7df3",
		00000245 => x"2b3a8ce8",
		00000246 => x"4230727a",
		00000247 => x"0f4df231",
		00000248 => x"50974f71",
		00000249 => x"1559c230",
		00000250 => x"66b1004c",
		00000251 => x"4b6e0548",
		00000252 => x"317083a2",
		00000253 => x"3751bf89",
		00000254 => x"07f17173",
		00000255 => x"5ee4e5f8",
		00000256 => x"1168f722",
		00000257 => x"3a34f078",
		00000258 => x"558fad04",
		00000259 => x"02a36cf3",
		00000260 => x"2cbdb767",
		00000261 => x"39908d4d",
		00000262 => x"6f7f753f",
		00000263 => x"5e855dd0",
		00000264 => x"5ebdb5ec",
		00000265 => x"5c2d6d94",
		00000266 => x"7d7f07a7",
		00000267 => x"5b02e86f",
		00000268 => x"559c5d3f",
		00000269 => x"39bf3df5",
		00000270 => x"26e31b9f",
		00000271 => x"36e9c262",
		00000272 => x"65431093",
		00000273 => x"631d0a1a",
		00000274 => x"039df59e",
		00000275 => x"144c43c6",
		00000276 => x"42c37c8f",
		00000277 => x"2994e447",
		00000278 => x"6f89dc42",
		00000279 => x"4227e5e7",
		00000280 => x"41e2511f",
		00000281 => x"473df528",
		00000282 => x"119563a6",
		00000283 => x"2bfa216a",
		00000284 => x"400403bb",
		00000285 => x"0d69599a",
		00000286 => x"45d18f29",
		00000287 => x"5cf84178",
		00000288 => x"2f3b68f0",
		00000289 => x"1cc9a9cf",
		00000290 => x"725c07ef",
		00000291 => x"48fbd534",
		00000292 => x"2b87c4f4",
		00000293 => x"0be2bc02",
		00000294 => x"22c8bfda",
		00000295 => x"77043528",
		00000296 => x"40ce7cbb",
		00000297 => x"1f2276f4",
		00000298 => x"1a04d186",
		00000299 => x"7178a854",
		00000300 => x"29392bd7",
		00000301 => x"21dcba7e",
		00000302 => x"32f73d92",
		00000303 => x"0581d526",
		00000304 => x"7818fc3e",
		00000305 => x"4011ef9c",
		00000306 => x"0a494bbd",
		00000307 => x"7a625ac5",
		00000308 => x"193a6792",
		00000309 => x"40a82208",
		00000310 => x"198931cb",
		00000311 => x"6109eaa6",
		00000312 => x"7f64d80b",
		00000313 => x"720e71a9",
		00000314 => x"72060509",
		00000315 => x"02324efb",
		00000316 => x"18da57c6",
		00000317 => x"22560269",
		00000318 => x"48459d85",
		00000319 => x"1d8f0cbb",
		00000320 => x"0ae48ec8",
		00000321 => x"4cd02369",
		00000322 => x"28946155",
		00000323 => x"0ab805b0",
		00000324 => x"2baa9d5a",
		00000325 => x"46fafe47",
		00000326 => x"44d2c38a",
		00000327 => x"11157793",
		00000328 => x"76f5bcd5",
		00000329 => x"71fc39d2",
		00000330 => x"678df2d4",
		00000331 => x"77bd07e3",
		00000332 => x"44601f4c",
		00000333 => x"11564b42",
		00000334 => x"649e4566",
		00000335 => x"737139e7",
		00000336 => x"3df25eaf",
		00000337 => x"3f034223",
		00000338 => x"5d830030",
		00000339 => x"32fd5553",
		00000340 => x"63733e4f",
		00000341 => x"039cdd0e",
		00000342 => x"20e0848c",
		00000343 => x"5b5c9813",
		00000344 => x"6a98702c",
		00000345 => x"6a034cba",
		00000346 => x"49fa131d",
		00000347 => x"6efed382",
		00000348 => x"3e392dc3",
		00000349 => x"2b96376d",
		00000350 => x"32aa02bb",
		00000351 => x"750e478c",
		00000352 => x"1cb0f0df",
		00000353 => x"6b9044a0",
		00000354 => x"4029351d",
		00000355 => x"76650e50",
		00000356 => x"10243fb4",
		00000357 => x"4e0c5128",
		00000358 => x"51408fb8",
		00000359 => x"00c35167",
		00000360 => x"72fa743f",
		00000361 => x"659adf17",
		00000362 => x"652ff4fd",
		00000363 => x"4cf40886",
		00000364 => x"4df8e1df",
		00000365 => x"7c3478c5",
		00000366 => x"3f4af01e",
		00000367 => x"2bf45a51",
		00000368 => x"590f63e5",
		00000369 => x"4ad4f423",
		00000370 => x"0fa80faf",
		00000371 => x"587b861d",
		00000372 => x"06b633cb",
		00000373 => x"2e29a37d",
		00000374 => x"6e4a7382",
		00000375 => x"3afa3b83",
		00000376 => x"2e50ceee",
		00000377 => x"7a955deb",
		00000378 => x"55a01097",
		00000379 => x"6d8ae2df",
		00000380 => x"35db84bf",
		00000381 => x"28628565",
		00000382 => x"2de8eab0",
		00000383 => x"1bb95cfc",
		00000384 => x"6298bb0c",
		00000385 => x"397a5dff",
		00000386 => x"2be883b0",
		00000387 => x"67ddef82",
		00000388 => x"6079b2f1",
		00000389 => x"18a2dc0b",
		00000390 => x"69056d5d",
		00000391 => x"7f9fc1df",
		00000392 => x"17206494",
		00000393 => x"30f1a5b7",
		00000394 => x"7d15e318",
		00000395 => x"672de6e0",
		00000396 => x"07fe1b0d",
		00000397 => x"6bba61f7",
		00000398 => x"3515c93a",
		00000399 => x"300afad7",
		00000400 => x"400f8ee7",
		00000401 => x"21fb3928",
		00000402 => x"6a2864ee",
		00000403 => x"7653a487",
		00000404 => x"16626ca6",
		00000405 => x"6d9c4528",
		00000406 => x"478e4f76",
		00000407 => x"302e0449",
		00000408 => x"2f2b924c",
		00000409 => x"08da35a7",
		00000410 => x"75f9b410",
		00000411 => x"25e004b5",
		00000412 => x"0fa86775",
		00000413 => x"74405021",
		00000414 => x"21f92756",
		00000415 => x"405cb83e",
		00000416 => x"68ef4a86",
		00000417 => x"4d7f6f41",
		00000418 => x"293ef6d2",
		00000419 => x"070757a9",
		00000420 => x"78dc3c46",
		00000421 => x"30b70347",
		00000422 => x"069af50a",
		00000423 => x"4b0107cb",
		00000424 => x"31b7afa5",
		00000425 => x"2635b5e7",
		00000426 => x"0dc1715d",
		00000427 => x"3b97149d",
		00000428 => x"49697108",
		00000429 => x"61ff05e1",
		00000430 => x"7b47aa8e",
		00000431 => x"5a69665f",
		00000432 => x"298f9c37",
		00000433 => x"1f0fe27b",
		00000434 => x"52cb8441",
		00000435 => x"39039e1a",
		00000436 => x"22097af3",
		00000437 => x"6ba0f64a",
		00000438 => x"38386a5e",
		00000439 => x"4808bb9e",
		00000440 => x"49279a87",
		00000441 => x"2c09f0e1",
		00000442 => x"1fcc01dd",
		00000443 => x"7971e50b",
		00000444 => x"586143a6",
		00000445 => x"3a4d5f24",
		00000446 => x"4020a179",
		00000447 => x"49983e0a",
		00000448 => x"73e637c8",
		00000449 => x"7625ba95",
		00000450 => x"2333e5a0",
		00000451 => x"2b28a8bc",
		00000452 => x"7a38ad31",
		00000453 => x"063e0cbe",
		00000454 => x"17528555",
		00000455 => x"0fc9959d",
		00000456 => x"028c7bd0",
		00000457 => x"36cca2b2",
		00000458 => x"5481961c",
		00000459 => x"3f8bf148",
		00000460 => x"5debee25",
		00000461 => x"10e1c065",
		00000462 => x"3d18e112",
		00000463 => x"447e57d8",
		00000464 => x"0579297e",
		00000465 => x"3c330d12",
		00000466 => x"7fc2dcc4",
		00000467 => x"455d6227",
		00000468 => x"121e5e39",
		00000469 => x"29b5289b",
		00000470 => x"6f6b789a",
		00000471 => x"2f54fb54",
		00000472 => x"721dbdbb",
		00000473 => x"788b253f",
		00000474 => x"1c450ad7",
		00000475 => x"4c811f19",
		00000476 => x"6e958dc9",
		00000477 => x"041d9d74",
		00000478 => x"3b50e5f5",
		00000479 => x"4086e1aa",
		00000480 => x"7325852c",
		00000481 => x"7460f3c8",
		00000482 => x"719a5dfc",
		00000483 => x"4cfa613e",
		00000484 => x"631c2db5",
		00000485 => x"79037121",
		00000486 => x"24f47506",
		00000487 => x"5a55faa8",
		00000488 => x"4a40dff4",
		00000489 => x"735130ac",
		00000490 => x"7d9baecb",
		00000491 => x"01c8b7c2",
		00000492 => x"290a2fb4",
		00000493 => x"5d6b89fb",
		00000494 => x"3178dc5b",
		00000495 => x"1d213ee5",
		00000496 => x"58100895",
		00000497 => x"71a0fd82",
		00000498 => x"080471d1",
		00000499 => x"6f902af5",
		00000500 => x"206e2a1c",
		00000501 => x"247de8c3",
		00000502 => x"1581b10d",
		00000503 => x"7f6a414e",
		00000504 => x"354158a5",
		00000505 => x"2dc6ada1",
		00000506 => x"3665a118",
		00000507 => x"058e56e9",
		00000508 => x"4db4183b",
		00000509 => x"01a902eb",
		00000510 => x"3f9775bf",
		00000511 => x"563e1734",
		00000512 => x"15172b17",
		00000513 => x"195ff47d",
		00000514 => x"05f7ade7",
		00000515 => x"227d54ad",
		00000516 => x"432bbc4c",
		00000517 => x"153d24f4",
		00000518 => x"61c60e48",
		00000519 => x"5e49a8b5",
		00000520 => x"76a4759c",
		00000521 => x"43ff6530",
		00000522 => x"6b7944c4",
		00000523 => x"18d6dd70",
		00000524 => x"26c09a9b",
		00000525 => x"3ffab6f9",
		00000526 => x"6ece6170",
		00000527 => x"70295d40",
		00000528 => x"3bd37c79",
		00000529 => x"1cb080f7",
		00000530 => x"2427396b",
		00000531 => x"438f4ae4",
		00000532 => x"0bcbdb7d",
		00000533 => x"0d36931e",
		00000534 => x"38aaccee",
		00000535 => x"4e723d6a",
		00000536 => x"45c14b3b",
		00000537 => x"4758fdf7",
		00000538 => x"23c014e4",
		00000539 => x"67580ca3",
		00000540 => x"18ff8d40",
		00000541 => x"42a68349",
		00000542 => x"786f1947",
		00000543 => x"76087696",
		00000544 => x"08acd93b",
		00000545 => x"5157abb8",
		00000546 => x"783e0168",
		00000547 => x"32399c0e",
		00000548 => x"340556fe",
		00000549 => x"661d475b",
		00000550 => x"6550747d",
		00000551 => x"396a4709",
		00000552 => x"0e338bbc",
		00000553 => x"07b30ebe",
		00000554 => x"48f602ad",
		00000555 => x"37616079",
		00000556 => x"617f430c",
		00000557 => x"53b92c10",
		00000558 => x"37cf3b7c",
		00000559 => x"42369b70",
		00000560 => x"2da0af9a",
		00000561 => x"13b1486b",
		00000562 => x"3f21cb44",
		00000563 => x"1139476b",
		00000564 => x"18e40ff8",
		00000565 => x"76fd7a3b",
		00000566 => x"1b16b18b",
		00000567 => x"7d0c809e",
		00000568 => x"1ee34bc5",
		00000569 => x"7c778620",
		00000570 => x"04cea81d",
		00000571 => x"1f4b172e",
		00000572 => x"747babb4",
		00000573 => x"1aa578dc",
		00000574 => x"09667ab6",
		00000575 => x"33aad36f",
		00000576 => x"76ac7640",
		00000577 => x"034f784d",
		00000578 => x"016702b6",
		00000579 => x"34c3ba22",
		00000580 => x"53fecd68",
		00000581 => x"2934a6d9",
		00000582 => x"4601b983",
		00000583 => x"03d565f1",
		00000584 => x"055b1195",
		00000585 => x"765ba802",
		00000586 => x"7881fbbf",
		00000587 => x"1f8e58ac",
		00000588 => x"5d89d8d3",
		00000589 => x"7181494f",
		00000590 => x"70875efa",
		00000591 => x"6d2bb7d2",
		00000592 => x"37c3d52f",
		00000593 => x"59731bec",
		00000594 => x"254c0b25",
		00000595 => x"76ad7129",
		00000596 => x"17cc7cb0",
		00000597 => x"26ef85b1",
		00000598 => x"0e6d97aa",
		00000599 => x"242a8839",
		00000600 => x"55e1af4a",
		00000601 => x"524ecb24",
		00000602 => x"6930a32c",
		00000603 => x"299381c4",
		00000604 => x"1b232e1f",
		00000605 => x"41fbbf0e",
		00000606 => x"0352dd08",
		00000607 => x"5fd434ff",
		00000608 => x"2e46b506",
		00000609 => x"649e2ad9",
		00000610 => x"139165b8",
		00000611 => x"3ba27676",
		00000612 => x"1ccaa2fa",
		00000613 => x"3507669a",
		00000614 => x"1c6c1fc4",
		00000615 => x"4159cf9a",
		00000616 => x"54ca398c",
		00000617 => x"75c45d64",
		00000618 => x"37a113f3",
		00000619 => x"320196b8",
		00000620 => x"47bdfce7",
		00000621 => x"182fc7ad",
		00000622 => x"31ee5d77",
		00000623 => x"09dd626a",
		00000624 => x"7de8ed07",
		00000625 => x"73baa8df",
		00000626 => x"3f9b8345",
		00000627 => x"6f290e8b",
		00000628 => x"0573bd75",
		00000629 => x"24b565b2",
		00000630 => x"11d20c48",
		00000631 => x"3ce1f481",
		00000632 => x"5d98a511",
		00000633 => x"5c383b36",
		00000634 => x"74d0f9b7",
		00000635 => x"0dacee22",
		00000636 => x"102012c5",
		00000637 => x"0f9dd73f",
		00000638 => x"3ae4b35a",
		00000639 => x"7696a08f",
		00000640 => x"6e5af5a5",
		00000641 => x"2d2b4aa9",
		00000642 => x"46a163a3",
		00000643 => x"4eab877d",
		00000644 => x"023ae71f",
		00000645 => x"38f6c8f8",
		00000646 => x"42abf130",
		00000647 => x"2d2f4df5",
		00000648 => x"24f5f9ce",
		00000649 => x"2e6fffb8",
		00000650 => x"1b4fd233",
		00000651 => x"31febac1",
		00000652 => x"77e31678",
		00000653 => x"060bcfcd",
		00000654 => x"0d8875e8",
		00000655 => x"41172f6c",
		00000656 => x"6a33a014",
		00000657 => x"714de6e9",
		00000658 => x"60629f99",
		00000659 => x"0c244400",
		00000660 => x"4be1a13e",
		00000661 => x"550c35f4",
		00000662 => x"299526bc",
		00000663 => x"5e39b833",
		00000664 => x"0a983900",
		00000665 => x"63e7c350",
		00000666 => x"559970fd",
		00000667 => x"1a5c9b0c",
		00000668 => x"7ac7e8cf",
		00000669 => x"3130335b",
		00000670 => x"170393aa",
		00000671 => x"359ae6cb",
		00000672 => x"10259574",
		00000673 => x"702bab8e",
		00000674 => x"3cd22deb",
		00000675 => x"11fe4752",
		00000676 => x"6cf9460a",
		00000677 => x"6e6f5be8",
		00000678 => x"00ae2bf8",
		00000679 => x"14cef667",
		00000680 => x"64f880a4",
		00000681 => x"65a27d67",
		00000682 => x"0b0c1852",
		00000683 => x"2a5f084e",
		00000684 => x"04221d6a",
		00000685 => x"0c923092",
		00000686 => x"12bd8942",
		00000687 => x"1c0a9506",
		00000688 => x"3a92d7e8",
		00000689 => x"3710f801",
		00000690 => x"77ee4e77",
		00000691 => x"19b480f3",
		00000692 => x"54a5a9ba",
		00000693 => x"33cc167b",
		00000694 => x"07a1ceb1",
		00000695 => x"07371ff9",
		00000696 => x"136ad299",
		00000697 => x"0ea4378f",
		00000698 => x"3b0d0300",
		00000699 => x"590c97ab",
		00000700 => x"0b8e8938",
		00000701 => x"1131b78b",
		00000702 => x"558c7aeb",
		00000703 => x"05455614",
		00000704 => x"2df18381",
		00000705 => x"3840b206",
		00000706 => x"7a60ba87",
		00000707 => x"67f03837",
		00000708 => x"68ebf276",
		00000709 => x"1a69a663",
		00000710 => x"68906a80",
		00000711 => x"1e9c3195",
		00000712 => x"1e18d6d9",
		00000713 => x"64738263",
		00000714 => x"3734ddc8",
		00000715 => x"2bb4dfe1",
		00000716 => x"55f687c0",
		00000717 => x"124e09a6",
		00000718 => x"0b718f42",
		00000719 => x"566f7f97",
		00000720 => x"0138a7ad",
		00000721 => x"2555f4f0",
		00000722 => x"29e7a6b5",
		00000723 => x"55a6da3e",
		00000724 => x"334a845e",
		00000725 => x"2c3b24d3",
		00000726 => x"64b8e34e",
		00000727 => x"1d4caea3",
		00000728 => x"684685fc",
		00000729 => x"07cac087",
		00000730 => x"076b12eb",
		00000731 => x"466bdb08",
		00000732 => x"0844e8dc",
		00000733 => x"0e1f3c00",
		00000734 => x"765f1cf0",
		00000735 => x"1ff566aa",
		00000736 => x"24df695e",
		00000737 => x"1e0337a6",
		00000738 => x"1003bfc5",
		00000739 => x"4756c633",
		00000740 => x"6574b1ae",
		00000741 => x"001a5cb2",
		00000742 => x"647a7cbe",
		00000743 => x"71441f61",
		00000744 => x"4d66997c",
		00000745 => x"728437ed",
		00000746 => x"623ad72e",
		00000747 => x"5206300e",
		00000748 => x"6e074c9a",
		00000749 => x"705c1572",
		00000750 => x"6d338b37",
		00000751 => x"45856f1a",
		00000752 => x"21b29687",
		00000753 => x"7544cf1b",
		00000754 => x"35df2275",
		00000755 => x"7cfe4240",
		00000756 => x"7e024c56",
		00000757 => x"471028e1",
		00000758 => x"2f124383",
		00000759 => x"2f702de0",
		00000760 => x"5023ac16",
		00000761 => x"10ac10df",
		00000762 => x"6c5a3701",
		00000763 => x"355bdf43",
		00000764 => x"703b54f5",
		00000765 => x"04409d91",
		00000766 => x"4d23c248",
		00000767 => x"2508ba63",
		00000768 => x"2cc80efc",
		00000769 => x"281fe6d6",
		00000770 => x"5859854d",
		00000771 => x"6bbb2a6e",
		00000772 => x"006bb17a",
		00000773 => x"6675df7f",
		00000774 => x"2cde9295",
		00000775 => x"40d07c03",
		00000776 => x"61220cb9",
		00000777 => x"005efd8e",
		00000778 => x"52c3ebd4",
		00000779 => x"25a636bc",
		00000780 => x"0a39ab53",
		00000781 => x"30736c11",
		00000782 => x"5c1c7c71",
		00000783 => x"17824676",
		00000784 => x"4e14ca18",
		00000785 => x"29ae8dc7",
		00000786 => x"38ec86a8",
		00000787 => x"6e17fcf0",
		00000788 => x"0d642127",
		00000789 => x"5de11a08",
		00000790 => x"4c54892d",
		00000791 => x"7a70a191",
		00000792 => x"5f6f0c09",
		00000793 => x"445bacdc",
		00000794 => x"196fd5ff",
		00000795 => x"3314c8e3",
		00000796 => x"514495c8",
		00000797 => x"56d521ab",
		00000798 => x"0909b2ec",
		00000799 => x"1888f755",
		00000800 => x"1a48aa0f",
		00000801 => x"5c743fbc",
		00000802 => x"2ddbb2d9",
		00000803 => x"36b41a62",
		00000804 => x"63962dc7",
		00000805 => x"3d8d0409",
		00000806 => x"2443291a",
		00000807 => x"53a55ba8",
		00000808 => x"71f5e0b3",
		00000809 => x"46c2fdf9",
		00000810 => x"7dd62717",
		00000811 => x"45b7f8b2",
		00000812 => x"14e8d6ef",
		00000813 => x"3192b2a4",
		00000814 => x"036b643c",
		00000815 => x"21539d3f",
		00000816 => x"5d46b849",
		00000817 => x"03fbaa49",
		00000818 => x"61d6f558",
		00000819 => x"74f5c737",
		00000820 => x"73516b84",
		00000821 => x"500c802d",
		00000822 => x"56135d50",
		00000823 => x"14a74c17",
		00000824 => x"63da4f36",
		00000825 => x"18a99693",
		00000826 => x"2ec95cdd",
		00000827 => x"178d6516",
		00000828 => x"0ce7737f",
		00000829 => x"1174fd9b",
		00000830 => x"7ffd2901",
		00000831 => x"5b73159c",
		00000832 => x"4d6696e8",
		00000833 => x"0cfa817a",
		00000834 => x"229e1de2",
		00000835 => x"0f854de3",
		00000836 => x"72460f94",
		00000837 => x"75073c16",
		00000838 => x"096b778f",
		00000839 => x"2e38dc6a",
		00000840 => x"074499ca",
		00000841 => x"7513caf4",
		00000842 => x"209ef5bf",
		00000843 => x"2e3a3803",
		00000844 => x"10a6d3e6",
		00000845 => x"2043e36f",
		00000846 => x"34936148",
		00000847 => x"0bdfc0eb",
		00000848 => x"4f7f7e23",
		00000849 => x"21471eaf",
		00000850 => x"427c56a0",
		00000851 => x"656e0a95",
		00000852 => x"46e02f9e",
		00000853 => x"6e9a5323",
		00000854 => x"0f47c754",
		00000855 => x"55470db6",
		00000856 => x"4478bd84",
		00000857 => x"0f7b663d",
		00000858 => x"7cd214c7",
		00000859 => x"754b5b63",
		00000860 => x"2a36898c",
		00000861 => x"24b918ff",
		00000862 => x"664dbd44",
		00000863 => x"668790e2",
		00000864 => x"51a98668",
		00000865 => x"6ee79b0c",
		00000866 => x"618b2a43",
		00000867 => x"7dd01ac3",
		00000868 => x"54379f7d",
		00000869 => x"277a0caa",
		00000870 => x"3841ca96",
		00000871 => x"7a76aa02",
		00000872 => x"1e13ba72",
		00000873 => x"00af5541",
		00000874 => x"0bfa11cd",
		00000875 => x"6b5e037b",
		00000876 => x"0e7ed276",
		00000877 => x"4f45cd96",
		00000878 => x"0ceb2660",
		00000879 => x"775571e9",
		00000880 => x"623885db",
		00000881 => x"3870d6c1",
		00000882 => x"6b2d152f",
		00000883 => x"31b26af0",
		00000884 => x"68a7ab47",
		00000885 => x"76d3ffe1",
		00000886 => x"71410885",
		00000887 => x"728c1400",
		00000888 => x"2dec2063",
		00000889 => x"78b37a0d",
		00000890 => x"5648851c",
		00000891 => x"1713e6ea",
		00000892 => x"68feeefb",
		00000893 => x"73c3921c",
		00000894 => x"10ef586c",
		00000895 => x"3196de1a",
		00000896 => x"000b6a9f",
		00000897 => x"352a7fdc",
		00000898 => x"1ad600b6",
		00000899 => x"1eb7be2f",
		00000900 => x"7537bffc",
		00000901 => x"008c0388",
		00000902 => x"6761d066",
		00000903 => x"3567129a",
		00000904 => x"10981ec6",
		00000905 => x"66c6cbc7",
		00000906 => x"6c703326",
		00000907 => x"0abbc6ed",
		00000908 => x"165afcf9",
		00000909 => x"449fd2d8",
		00000910 => x"2222a1d2",
		00000911 => x"35ed3e26",
		00000912 => x"1585dfe9",
		00000913 => x"63819691",
		00000914 => x"7124ef48",
		00000915 => x"31efdcd9",
		00000916 => x"69fe1e67",
		00000917 => x"271d1bff",
		00000918 => x"084f401d",
		00000919 => x"6fd5a302",
		00000920 => x"030cc671",
		00000921 => x"0f9e37dd",
		00000922 => x"65472564",
		00000923 => x"48d3985f",
		00000924 => x"326463fb",
		00000925 => x"22100730",
		00000926 => x"48c213ff",
		00000927 => x"06db0ff5",
		00000928 => x"51ad94c4",
		00000929 => x"565e5448",
		00000930 => x"459498ea",
		00000931 => x"5b6e98c8",
		00000932 => x"18103ba3",
		00000933 => x"7000e32f",
		00000934 => x"27b8f977",
		00000935 => x"27dc26f2",
		00000936 => x"4c791fd2",
		00000937 => x"46114fe4",
		00000938 => x"64637e75",
		00000939 => x"54b63a2e",
		00000940 => x"2b4abaf3",
		00000941 => x"7f1cc6ac",
		00000942 => x"02e68cfd",
		00000943 => x"5531cda9",
		00000944 => x"129817dd",
		00000945 => x"2770475e",
		00000946 => x"24771c9a",
		00000947 => x"70ab2695",
		00000948 => x"7b07baf8",
		00000949 => x"19986d75",
		00000950 => x"36a72531",
		00000951 => x"1b21be74",
		00000952 => x"3fade224",
		00000953 => x"05c178cf",
		00000954 => x"361bc1d4",
		00000955 => x"08679efe",
		00000956 => x"6edc69a9",
		00000957 => x"664ace47",
		00000958 => x"667b35d5",
		00000959 => x"7c569375",
		00000960 => x"13b4dfdf",
		00000961 => x"15c79bbe",
		00000962 => x"5541e2f1",
		00000963 => x"060f5663",
		00000964 => x"4662750a",
		00000965 => x"1c76d682",
		00000966 => x"72e1bc3c",
		00000967 => x"6a2625bf",
		00000968 => x"0807918c",
		00000969 => x"3978090b",
		00000970 => x"4a056bcf",
		00000971 => x"7b8817a1",
		00000972 => x"184c01bb",
		00000973 => x"334ac03a",
		00000974 => x"48e043b4",
		00000975 => x"5bf296fe",
		00000976 => x"68992c61",
		00000977 => x"6e4e9da3",
		00000978 => x"378e32b8",
		00000979 => x"5b06ab94",
		00000980 => x"447448c2",
		00000981 => x"782eac59",
		00000982 => x"2ebc801f",
		00000983 => x"098caf11",
		00000984 => x"78f05861",
		00000985 => x"6a5c088b",
		00000986 => x"6e63741d",
		00000987 => x"1bac0541",
		00000988 => x"0b7afd6a",
		00000989 => x"383b957b",
		00000990 => x"05783bb9",
		00000991 => x"782eae07",
		00000992 => x"4478b0f0",
		00000993 => x"76813066",
		00000994 => x"27dde237",
		00000995 => x"59c46888",
		00000996 => x"03ff8495",
		00000997 => x"1aa75f7e",
		00000998 => x"566d31c5",
		00000999 => x"048fb6fa",
		00001000 => x"13fde11a",
		00001001 => x"6d7ad467",
		00001002 => x"5268d0b7",
		00001003 => x"433de2ba",
		00001004 => x"0c9f4de4",
		00001005 => x"7d35224c",
		00001006 => x"5b61ea20",
		00001007 => x"067f5317",
		00001008 => x"6b3191f5",
		00001009 => x"34b54afa",
		00001010 => x"6609bd6e",
		00001011 => x"5d995bc8",
		00001012 => x"71049498",
		00001013 => x"3c7ad0a7",
		00001014 => x"4ec0ff7d",
		00001015 => x"3131f218",
		00001016 => x"2ab89b7f",
		00001017 => x"54b96778",
		00001018 => x"175a350a",
		00001019 => x"524b443d",
		00001020 => x"5434832b",
		00001021 => x"33cd592c",
		00001022 => x"7cb49421",
		00001023 => x"36dd81d8"
	);

end package neorv32_dcache_memory_tb_pkg;
